`ifndef _{{name.upper()}}_TYPES_SVH_
    `define _{{name.upper()}}_TYPES_SVH_

    typedef virtual /*interface*/ virtual_interface;

`endif