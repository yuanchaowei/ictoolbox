module xmpl_dsp_msf #(
)(
    // 123
    input                           clk_i,
    input                           reset_n_i,

    // wd1
    input                           xmpl_dsp_msf_a_i,
    input  [12 - 1 : 0]             xmpl_dsp_msf_b_i, //asdwad

    // 1df1234
    input  [32 - 1 : 0]             xmpl_dsp_msf_c_o,
    input  [32 - 1 : 0]             xmpl_dsp_msf_status_o

);

logic [32 - 1 : 0] sadwd;
logic              sxawd;
logic              123;
//awudhiuwha
