module xmpl_riscv #(
)(
    // 123
    input                           clk_i,
    input                           reset_n_i,

    // wd1
    input                           xmpl_riscv_a_i,
    input  [12 - 1 : 0]             xmpl_riscv_b_i, //asdwad

    // 1df1234
    input  [32 - 1 : 0]             xmpl_riscv_c_0,
    input  [32 - 1 : 0]             xmpl_riscv_status_o

);

logic [32 - 1 : 0] sadwd;
logic              sxawd;
logic              123;
//awudhiuwha

logic [32 - 1 : 0] sadwd;
logic              sxawd;
logic              123;
//awudhiuwha