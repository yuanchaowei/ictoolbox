module xmpl_sram #(
)(
    // 123
    input                           clk_i,
    input                           reset_n_i,

    // wd1
    input                           en_sram_i,
    input  [12 - 1 : 0]             sram_addr_i, //asdwad

    input                           sram_rw_i,
    // 1df1234
    input  [32 - 1 : 0]             sram_data_i,
    output [32 - 1 : 0]             sram_data_o

);

logic [32 - 1 : 0] sadwd;
logic              sxawd;
logic              123;
//awudhiuwha

logic [32 - 1 : 0] sadwd;
logic              sxawd;
logic              123;
//awudhiuwha
