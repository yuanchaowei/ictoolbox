module xmpl_loongson #(
)(
    input  [32 - 1 : 0] xmpl_loongson_i,
    input  [32 - 1 : 0] xmpl_stone2loongson_i,
    output [32 - 1 : 0] xmpl_loongson2stone_o

);

logic [32 - 1 : 0] sadwd;
logic              sxawd;
logic              123;
//awudhiuwha
