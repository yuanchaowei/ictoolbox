`ifndef _{{name.upper()}}_DEF_SVH_
	`define _{{name.upper()}}_DEF_SVH_

    
    
`endif