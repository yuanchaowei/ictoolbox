module xmpl_stone #(
)(
    input  [32 - 1 : 0] xmpl_stone_i,
    input  [32 - 1 : 0] xmpl_loongson2stone_i,
    output [32 - 1 : 0] xmpl_stone2loongson_o
);

logic [32 - 1 : 0] sadwd;
logic              sxawd;
logic              123;
//awudhiuwha

logic [32 - 1 : 0] sadwd;
logic              sxawd;
logic              123;
//awudhiuwha
