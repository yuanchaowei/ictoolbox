module xmpl_clkgating #(
)(
    input a_i,
    input en_i,
    output c_o
)
